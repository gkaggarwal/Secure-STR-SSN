----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06.12.2024 19:33:10
-- Design Name: 
-- Module Name: Design_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Design_tb is
    -- No ports for the testbench
--    generic (
--    pattern :  std_logic_vector(129 downto 0):=(others=>'0')
--  );
  
end Design_tb;

architecture Behavioral of Design_tb is

    -- Generic parameter for 16 key the pattern

constant key_size : integer := 16;
    --signal pattern : std_logic_vector(key_size + 1 downto 0):="010110100100001101111011110111111010011100111110110101100110111001111101010101000111101010100011011010111101111011111100010111000011000010000110001111010101111100010100110011011101001000110101010010011001101111000101101001100001110001111111010111111111111101";
    signal data : std_logic_vector(key_size - 1 downto 0):="0010001011011101";
    
    --signal pattern2 : std_logic_vector(key_size + 1 downto 0):= "010110011100001110010110110100010000101010110110001101101010001100000001110111011101110011000111010010110011110111110100100101110001011010010000111011010010011100111101110111011111010000011111110111011100001000101001001001101010101111111000111111000001100011";
   -- signal pattern3 : std_logic_vector(key_size + 1 downto 0):= "011010110111111110110100000010001101000111101100100100000010011001111001001001000110100000001100100111001100100111001011110010101010001001010111100000001101100000100110111101100100111110101100100111001100101100101101011000000111001111001101000101100000101001";
    --signal pattern4 : std_logic_vector(key_size + 1 downto 0):= "011000001111101001000011000011101010110001001110010010001001000011101001011101011000010111000100001011011010001100100010011010101011110001001110110001011010001101100000000101011010010111001111001101001111111010101101111111000000011110111000110111101111111100";
    --signal pattern5 : std_logic_vector(key_size + 1 downto 0):= "011010001001000001111000100101110010111100100111111100100111000101110001010100101110100101001110000110010011100011010110011011110010000101010011101100010110000000100101000000001110101001001010100010110011111011010111011010000011001100101111111100101110010101";
   -- signal pattern6 : std_logic_vector(key_size + 1 downto 0):= "011111011010100111011100111010111110000001100000010010110011001111111101010001100111011010010101000001011100011111110010010011000101111011010011010111100110000111101101101111110101011110110001110001110010010101100011000111011010110000011001001011100010011001";
  --  signal pattern : std_logic_vector(key_size + 1 downto 0):= "011101001100100100000111000000000110000110001101101111000101011100001000110111010100001011101000011111111010101110001100111100010110110010100011000011011111101100001001010100011110101010011110111110011111001110101100101000101101110100110011110000001100000110";
   --  signal pattern : std_logic_vector(key_size + 1 downto 0):= "011001000010001101011010100001101110111001011001100000100011000000101010111010111101100111111010100110010000111011110011010110001001001010100110011101010001101101010110010111101101111101011100110110100110111000110011101010011100010010110011111110010111111101";
   -- signal pattern : std_logic_vector(key_size + 1 downto 0):= "011111001011111101000100110001100111101110101010000101010001111001110010011101010111111101100100010111001100110001101100100011001001111011101010011000000001101011100100110000011001011101000011101111010100010011111110110011010111000100110110111010110110100010";
    signal pattern : std_logic_vector(key_size + 1 downto 0):= "010010001110010111";
    
 
 
 
    -- Signals to connect to the DUT (Device Under Test)
    signal TCLK, TMS, TDI, TDO : std_logic;
    constant CLK_PERIOD : time := 100 ns;

    -- Instantiate the Design Under Test (DUT)
    component Design is
        generic (
            key_size : integer := 4;
            Data :STD_LOGIC_VECTOR := "1010";
            seed_value : std_logic_vector := "0101" -- Generic seed value
        );
        port (
            TCLK, TMS, TDI : in std_logic;
            TDO : out std_logic
        );
    end component;
--seed 1 1100000000000011110000001001001000101011101110010001101010101101111111010011011100110101010111100100001111110001001010001100010100010011100100000110001100011110110100111111100010011111111100001010011010101111011000010100101110000011000110001101000110111011
--seed 2 0100101000010000010010000001111111101011011011110011000100110011000000100001110000110011001100010100101101110110010001101110111001001110110111000011000101011101110010010101001100110011001000000101001111101101001011011111110001100111011011101001000100101010
--seed 3 1011110000101110011101010001010010000010111101110101110101010010110101111000010110101100011010110000101101000000100011111011001111111101000111010010110101010010110101000000111010011011011010001010101100000110110101100010011101001100000111011000000011011110
--seed 4 0100000001100011010010011000100000010000001101111110000001011101010001010011101110111110000000101101001110111001011001011001000111111110101100110101001110110111000110010011100010111100111011100100011011001101101001011001011111100100010100011011100001000011
--seed 5 1111101001110100000001110101010100001110110011110110000101011100111111011011111001000000011110110000001011100101100101111110001101000110101011110100100101101010001001011110111001110111111001001110010010110100000010110100011101001110110010001000011011001110
--seed 6 1010101100100111011010100001011110110010010100101111101101001001001001011000111111000001101101100010001010100011110101110110001110010101101101000000100100111000011111101110110010101001111100000001010101011101100000101000001000011110010100110010111110110000
--seed 7 1010000101000001000101010111001101110011110101111001010000101000011000101111111000100111111011000101100000110100010100111101011011100100010101001001111110000000100011100111000111110011010011000100111110010001101101001010001010000000010010000110110101011100
--seed 8 1100000011101000000101011101100100101111100101010010011010111011010100111100001101100011101011111101101001111100101010111111011011001011110101000110010001101010111110000010101100011110011111110000010100110000101010111010011001101000111110111101001100011010
--seed 9 1100111011011110011011010110010011110101011000000101100111110001100100011100111010100001010110100111101000000010101111100110001011010100110101101001010101010011100110101100000011111100101101001010001001111110001111111001100010101001010110011100000111010000
--seed 10 1011101001001111011001101011011101101110110110010001011000001000110100100001101001101101001100100110010100101110001100100001010110000100011000111111000001101001110111101000111111011000110011101010101011000000100010010010001010000110110011000100011011001100




begin
    -- Instantiate the DUT
    DUT: Design
        generic map (
            key_size => key_size,
            Data => data,
            seed_value => "0011101001001100"
        )
        port map (
            TCLK => TCLK,
            TMS  => TMS,
            TDI  => TDI,
            TDO  => TDO
        );

    -- Clock generation process
    clk_gen: process
    begin
        TCLK <= '0';
        wait for CLK_PERIOD / 2;
        TCLK <= '1';
        wait for CLK_PERIOD / 2;
    end process;

    -- Stimulus process
    stim_proc: process
        variable index : integer := key_size + 1; -- Start from MSB
    begin
        -- Apply reset
        TMS <= '0';
        TDI <= '0';
        wait for CLK_PERIOD;

        -- Test 1: Apply matching input bits
        TDI <= '1';
        TMS <= '1';
        wait for CLK_PERIOD;

        -- Apply the pattern
        while index >= 0 loop
            TDI <= pattern(index);
            TMS <= '0';
            wait for CLK_PERIOD; -- Apply on rising edge of clock
            index := index - 1;
        end loop;

        -- Perform additional operations if needed
  --- NOW DATA FOR UPDATE
           for i in 1 to 4 loop
        TDI <= '1';
        TMS <= '0';
        wait for CLK_PERIOD;

        TDI <= '1';
        TMS <= '0';
        wait for CLK_PERIOD;

        TDI <= '1';
        TMS <= '0';
        wait for CLK_PERIOD;

        TDI <= '1';
        TMS <= '0';
        wait for CLK_PERIOD;
    end loop;
    
--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;
--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;
--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;
--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;
        
        
        
        -- fOR UPDATE
        TDI <= '0';
        TMS <= '1';
        wait for CLK_PERIOD;
        
        TDI <= '0';
        TMS <= '1';
        wait for CLK_PERIOD;
        -- End simulation
    end process;

end Behavioral;


--    -- Generic parameter for 32 key the pattern

--constant key_size : integer := 32;
--    --signal pattern : std_logic_vector(key_size + 1 downto 0):="010110100100001101111011110111111010011100111110110101100110111001111101010101000111101010100011011010111101111011111100010111000011000010000110001111010101111100010100110011011101001000110101010010011001101111000101101001100001110001111111010111111111111101";
--    signal data : std_logic_vector(key_size - 1 downto 0):="01001101101001111100100111000110";
    
--    --signal pattern2 : std_logic_vector(key_size + 1 downto 0):= "010110011100001110010110110100010000101010110110001101101010001100000001110111011101110011000111010010110011110111110100100101110001011010010000111011010010011100111101110111011111010000011111110111011100001000101001001001101010101111111000111111000001100011";
--   -- signal pattern3 : std_logic_vector(key_size + 1 downto 0):= "011010110111111110110100000010001101000111101100100100000010011001111001001001000110100000001100100111001100100111001011110010101010001001010111100000001101100000100110111101100100111110101100100111001100101100101101011000000111001111001101000101100000101001";
--    --signal pattern4 : std_logic_vector(key_size + 1 downto 0):= "011000001111101001000011000011101010110001001110010010001001000011101001011101011000010111000100001011011010001100100010011010101011110001001110110001011010001101100000000101011010010111001111001101001111111010101101111111000000011110111000110111101111111100";
--    --signal pattern5 : std_logic_vector(key_size + 1 downto 0):= "011010001001000001111000100101110010111100100111111100100111000101110001010100101110100101001110000110010011100011010110011011110010000101010011101100010110000000100101000000001110101001001010100010110011111011010111011010000011001100101111111100101110010101";
--   -- signal pattern6 : std_logic_vector(key_size + 1 downto 0):= "011111011010100111011100111010111110000001100000010010110011001111111101010001100111011010010101000001011100011111110010010011000101111011010011010111100110000111101101101111110101011110110001110001110010010101100011000111011010110000011001001011100010011001";
--  --  signal pattern : std_logic_vector(key_size + 1 downto 0):= "011101001100100100000111000000000110000110001101101111000101011100001000110111010100001011101000011111111010101110001100111100010110110010100011000011011111101100001001010100011110101010011110111110011111001110101100101000101101110100110011110000001100000110";
--   --  signal pattern : std_logic_vector(key_size + 1 downto 0):= "011001000010001101011010100001101110111001011001100000100011000000101010111010111101100111111010100110010000111011110011010110001001001010100110011101010001101101010110010111101101111101011100110110100110111000110011101010011100010010110011111110010111111101";
--   -- signal pattern : std_logic_vector(key_size + 1 downto 0):= "011111001011111101000100110001100111101110101010000101010001111001110010011101010111111101100100010111001100110001101100100011001001111011101010011000000001101011100100110000011001011101000011101111010100010011111110110011010111000100110110111010110110100010";
--    signal pattern : std_logic_vector(key_size + 1 downto 0):= "0111110000010110111011100001000010";
    
 
 
 
--    -- Signals to connect to the DUT (Device Under Test)
--    signal TCLK, TMS, TDI, TDO : std_logic;
--    constant CLK_PERIOD : time := 100 ns;

--    -- Instantiate the Design Under Test (DUT)
--    component Design is
--        generic (
--            key_size : integer := 4;
--            Data :STD_LOGIC_VECTOR := "1010";
--            seed_value : std_logic_vector := "0101" -- Generic seed value
--        );
--        port (
--            TCLK, TMS, TDI : in std_logic;
--            TDO : out std_logic
--        );
--    end component;
----seed 1 1100000000000011110000001001001000101011101110010001101010101101111111010011011100110101010111100100001111110001001010001100010100010011100100000110001100011110110100111111100010011111111100001010011010101111011000010100101110000011000110001101000110111011
----seed 2 0100101000010000010010000001111111101011011011110011000100110011000000100001110000110011001100010100101101110110010001101110111001001110110111000011000101011101110010010101001100110011001000000101001111101101001011011111110001100111011011101001000100101010
----seed 3 1011110000101110011101010001010010000010111101110101110101010010110101111000010110101100011010110000101101000000100011111011001111111101000111010010110101010010110101000000111010011011011010001010101100000110110101100010011101001100000111011000000011011110
----seed 4 0100000001100011010010011000100000010000001101111110000001011101010001010011101110111110000000101101001110111001011001011001000111111110101100110101001110110111000110010011100010111100111011100100011011001101101001011001011111100100010100011011100001000011
----seed 5 1111101001110100000001110101010100001110110011110110000101011100111111011011111001000000011110110000001011100101100101111110001101000110101011110100100101101010001001011110111001110111111001001110010010110100000010110100011101001110110010001000011011001110
----seed 6 1010101100100111011010100001011110110010010100101111101101001001001001011000111111000001101101100010001010100011110101110110001110010101101101000000100100111000011111101110110010101001111100000001010101011101100000101000001000011110010100110010111110110000
----seed 7 1010000101000001000101010111001101110011110101111001010000101000011000101111111000100111111011000101100000110100010100111101011011100100010101001001111110000000100011100111000111110011010011000100111110010001101101001010001010000000010010000110110101011100
----seed 8 1100000011101000000101011101100100101111100101010010011010111011010100111100001101100011101011111101101001111100101010111111011011001011110101000110010001101010111110000010101100011110011111110000010100110000101010111010011001101000111110111101001100011010
----seed 9 1100111011011110011011010110010011110101011000000101100111110001100100011100111010100001010110100111101000000010101111100110001011010100110101101001010101010011100110101100000011111100101101001010001001111110001111111001100010101001010110011100000111010000
----seed 10 1011101001001111011001101011011101101110110110010001011000001000110100100001101001101101001100100110010100101110001100100001010110000100011000111111000001101001110111101000111111011000110011101010101011000000100010010010001010000110110011000100011011001100




--begin
--    -- Instantiate the DUT
--    DUT: Design
--        generic map (
--            key_size => key_size,
--            Data => data,
--            seed_value => "11000110001001100110111000010000"
--        )
--        port map (
--            TCLK => TCLK,
--            TMS  => TMS,
--            TDI  => TDI,
--            TDO  => TDO
--        );

--    -- Clock generation process
--    clk_gen: process
--    begin
--        TCLK <= '0';
--        wait for CLK_PERIOD / 2;
--        TCLK <= '1';
--        wait for CLK_PERIOD / 2;
--    end process;

--    -- Stimulus process
--    stim_proc: process
--        variable index : integer := key_size + 1; -- Start from MSB
--    begin
--        -- Apply reset
--        TMS <= '0';
--        TDI <= '0';
--        wait for CLK_PERIOD;

--        -- Test 1: Apply matching input bits
--        TDI <= '1';
--        TMS <= '1';
--        wait for CLK_PERIOD;

--        -- Apply the pattern
--        while index >= 0 loop
--            TDI <= pattern(index);
--            TMS <= '0';
--            wait for CLK_PERIOD; -- Apply on rising edge of clock
--            index := index - 1;
--        end loop;

--        -- Perform additional operations if needed
--  --- NOW DATA FOR UPDATE
--           for i in 1 to 8 loop
--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;

--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;

--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;

--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;
--    end loop;
    
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
        
        
        
--        -- fOR UPDATE
--        TDI <= '0';
--        TMS <= '1';
--        wait for CLK_PERIOD;
        
--        TDI <= '0';
--        TMS <= '1';
--        wait for CLK_PERIOD;
--        -- End simulation
--    end process;

--end Behavioral;








    -- Generic parameter for 256 key the pattern
--    constant key_size : integer := 256;
--    --signal pattern : std_logic_vector(key_size + 1 downto 0):="010110100100001101111011110111111010011100111110110101100110111001111101010101000111101010100011011010111101111011111100010111000011000010000110001111010101111100010100110011011101001000110101010010011001101111000101101001100001110001111111010111111111111101";
--    signal data : std_logic_vector(key_size - 1 downto 0):="1010101010101010100101111010001100001000011110000100000000000010111001000011001000010110111111011000000100010001100110010001001001001010100000010100011100001110100101110100010110001010100000010010001001001100100111101111000010010011111100101001010110110000";
    
--    --signal pattern2 : std_logic_vector(key_size + 1 downto 0):= "010110011100001110010110110100010000101010110110001101101010001100000001110111011101110011000111010010110011110111110100100101110001011010010000111011010010011100111101110111011111010000011111110111011100001000101001001001101010101111111000111111000001100011";
--   -- signal pattern3 : std_logic_vector(key_size + 1 downto 0):= "011010110111111110110100000010001101000111101100100100000010011001111001001001000110100000001100100111001100100111001011110010101010001001010111100000001101100000100110111101100100111110101100100111001100101100101101011000000111001111001101000101100000101001";
--    --signal pattern4 : std_logic_vector(key_size + 1 downto 0):= "011000001111101001000011000011101010110001001110010010001001000011101001011101011000010111000100001011011010001100100010011010101011110001001110110001011010001101100000000101011010010111001111001101001111111010101101111111000000011110111000110111101111111100";
--    --signal pattern5 : std_logic_vector(key_size + 1 downto 0):= "011010001001000001111000100101110010111100100111111100100111000101110001010100101110100101001110000110010011100011010110011011110010000101010011101100010110000000100101000000001110101001001010100010110011111011010111011010000011001100101111111100101110010101";
--   -- signal pattern6 : std_logic_vector(key_size + 1 downto 0):= "011111011010100111011100111010111110000001100000010010110011001111111101010001100111011010010101000001011100011111110010010011000101111011010011010111100110000111101101101111110101011110110001110001110010010101100011000111011010110000011001001011100010011001";
--  --  signal pattern : std_logic_vector(key_size + 1 downto 0):= "011101001100100100000111000000000110000110001101101111000101011100001000110111010100001011101000011111111010101110001100111100010110110010100011000011011111101100001001010100011110101010011110111110011111001110101100101000101101110100110011110000001100000110";
--   --  signal pattern : std_logic_vector(key_size + 1 downto 0):= "011001000010001101011010100001101110111001011001100000100011000000101010111010111101100111111010100110010000111011110011010110001001001010100110011101010001101101010110010111101101111101011100110110100110111000110011101010011100010010110011111110010111111101";
--   -- signal pattern : std_logic_vector(key_size + 1 downto 0):= "011111001011111101000100110001100111101110101010000101010001111001110010011101010111111101100100010111001100110001101100100011001001111011101010011000000001101011100100110000011001011101000011101111010100010011111110110011010111000100110110111010110110100010";
--    signal pattern : std_logic_vector(key_size + 1 downto 0):= "011101110110111100001000100100000110000111000111100000001001100110010111011110110101011110010100101110010000001010100001000011111011001111100010000101100011000100011101110010010001101111100011011110000001001111000100100101101101001001101110110101110001101001";
    
 
 
 
--    -- Signals to connect to the DUT (Device Under Test)
--    signal TCLK, TMS, TDI, TDO : std_logic;
--    constant CLK_PERIOD : time := 100 ns;

--    -- Instantiate the Design Under Test (DUT)
--    component Design is
--        generic (
--            key_size : integer := 4;
--            Data :STD_LOGIC_VECTOR := "1010";
--            seed_value : std_logic_vector := "0101" -- Generic seed value
--        );
--        port (
--            TCLK, TMS, TDI : in std_logic;
--            TDO : out std_logic
--        );
--    end component;
----seed 1 1100000000000011110000001001001000101011101110010001101010101101111111010011011100110101010111100100001111110001001010001100010100010011100100000110001100011110110100111111100010011111111100001010011010101111011000010100101110000011000110001101000110111011
----seed 2 0100101000010000010010000001111111101011011011110011000100110011000000100001110000110011001100010100101101110110010001101110111001001110110111000011000101011101110010010101001100110011001000000101001111101101001011011111110001100111011011101001000100101010
----seed 3 1011110000101110011101010001010010000010111101110101110101010010110101111000010110101100011010110000101101000000100011111011001111111101000111010010110101010010110101000000111010011011011010001010101100000110110101100010011101001100000111011000000011011110
----seed 4 0100000001100011010010011000100000010000001101111110000001011101010001010011101110111110000000101101001110111001011001011001000111111110101100110101001110110111000110010011100010111100111011100100011011001101101001011001011111100100010100011011100001000011
----seed 5 1111101001110100000001110101010100001110110011110110000101011100111111011011111001000000011110110000001011100101100101111110001101000110101011110100100101101010001001011110111001110111111001001110010010110100000010110100011101001110110010001000011011001110
----seed 6 1010101100100111011010100001011110110010010100101111101101001001001001011000111111000001101101100010001010100011110101110110001110010101101101000000100100111000011111101110110010101001111100000001010101011101100000101000001000011110010100110010111110110000
----seed 7 1010000101000001000101010111001101110011110101111001010000101000011000101111111000100111111011000101100000110100010100111101011011100100010101001001111110000000100011100111000111110011010011000100111110010001101101001010001010000000010010000110110101011100
----seed 8 1100000011101000000101011101100100101111100101010010011010111011010100111100001101100011101011111101101001111100101010111111011011001011110101000110010001101010111110000010101100011110011111110000010100110000101010111010011001101000111110111101001100011010
----seed 9 1100111011011110011011010110010011110101011000000101100111110001100100011100111010100001010110100111101000000010101111100110001011010100110101101001010101010011100110101100000011111100101101001010001001111110001111111001100010101001010110011100000111010000
----seed 10 1011101001001111011001101011011101101110110110010001011000001000110100100001101001101101001100100110010100101110001100100001010110000100011000111111000001101001110111101000111111011000110011101010101011000000100010010010001010000110110011000100011011001100




--begin
--    -- Instantiate the DUT
--    DUT: Design
--        generic map (
--            key_size => key_size,
--            Data => data,
--            seed_value => "1011101001001111011001101011011101101110110110010001011000001000110100100001101001101101001100100110010100101110001100100001010110000100011000111111000001101001110111101000111111011000110011101010101011000000100010010010001010000110110011000100011011001100"
--        )
--        port map (
--            TCLK => TCLK,
--            TMS  => TMS,
--            TDI  => TDI,
--            TDO  => TDO
--        );

--    -- Clock generation process
--    clk_gen: process
--    begin
--        TCLK <= '0';
--        wait for CLK_PERIOD / 2;
--        TCLK <= '1';
--        wait for CLK_PERIOD / 2;
--    end process;

--    -- Stimulus process
--    stim_proc: process
--        variable index : integer := key_size + 1; -- Start from MSB
--    begin
--        -- Apply reset
--        TMS <= '0';
--        TDI <= '0';
--        wait for CLK_PERIOD;

--        -- Test 1: Apply matching input bits
--        TDI <= '1';
--        TMS <= '1';
--        wait for CLK_PERIOD;

--        -- Apply the pattern
--        while index >= 0 loop
--            TDI <= pattern(index);
--            TMS <= '0';
--            wait for CLK_PERIOD; -- Apply on rising edge of clock
--            index := index - 1;
--        end loop;

--        -- Perform additional operations if needed
--  --- NOW DATA FOR UPDATE
--           for i in 1 to 64 loop
--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;

--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;

--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;

--        TDI <= '1';
--        TMS <= '0';
--        wait for CLK_PERIOD;
--    end loop;
    
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
----        TDI <= '1';
----        TMS <= '0';
----        wait for CLK_PERIOD;
        
        
        
--        -- fOR UPDATE
--        TDI <= '0';
--        TMS <= '1';
--        wait for CLK_PERIOD;
        
--        TDI <= '0';
--        TMS <= '1';
--        wait for CLK_PERIOD;
--        -- End simulation
--    end process;

--end Behavioral;